module Slave_1 #(
  parameter                     ADD_WIDTH = 9,
  parameter                     WIDTH = 32
)(
  //Global Signals
  //---------------------------------------------------------------------------
  input                         Pclk,
  input                         Presetn,
  //---------------------------------------------------------------------------

  //From Master
  //---------------------------------------------------------------------------
  input                         Psel,
  input                         Penable,
  input                         Pwrite,
  input [ADD_WIDTH - 2 : 0]     Paddr,
  input [WIDTH - 1 : 0]         Pwdata,
  //---------------------------------------------------------------------------

  //To Master
  //---------------------------------------------------------------------------
  output reg [WIDTH - 1 : 0]    Prdata,
  output  Pready
  //---------------------------------------------------------------------------
);

  //Memory Depth calculation
  //---------------------------------------------------------------------------
  localparam DEPTH = 2 ** (ADD_WIDTH - 1);
  //---------------------------------------------------------------------------

  //Memory Definition
  //---------------------------------------------------------------------------
  reg [WIDTH - 1 : 0] mem [0 : DEPTH - 1];
  //---------------------------------------------------------------------------

  //Read Opration
  //---------------------------------------------------------------------------
  always @(posedge Pclk) begin
    if(!Presetn)
      Prdata <= 'b0;
    else begin
          if(Psel && Penable) begin
            if(!Pwrite)
          Prdata <=  mem[Paddr];
          end
          else begin
            Prdata <= 1'b0;
          end
    end
  end
  //---------------------------------------------------------------------------

  //write opertion
  //---------------------------------------------------------------------------
  always @(posedge Pclk) begin
    if(Psel && Penable) begin
            if(Pwrite)
          mem[Paddr] <= Pwdata;
          end
  end
  //---------------------------------------------------------------------------

  //Pready assignment based on sel and enable
  //---------------------------------------------------------------------------
  assign Pready = Psel && Penable;
  //---------------------------------------------------------------------------

endmodule
